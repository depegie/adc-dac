`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/25/2022 10:01:52 PM
// Design Name: 
// Module Name: Serializer_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Serializer_tb;

    logic Clk_tb;
    logic Rst_tb;
    logic [11 : 0] DATAIN_tb;
    logic SCLK_tb;
    logic SYNCn_tb;
    logic DIN_tb;
    
    Serializer serial(
        .Clk(Clk_tb),
        .Rst(Rst_tb),
        .DATAIN(DATAIN_tb),
        .SCLK(SCLK_tb),
        .SYNCn(SYNCn_tb),
        .DIN(DIN_tb)
    );
    
    always #4 Clk_tb = ~Clk_tb;
    
    initial begin
        Clk_tb = 0;
        Rst_tb = 0;
        DATAIN_tb = 12'b1100_1001_0011;
        #5000 DATAIN_tb = 12'b1000_1001_0101;
        #5000 DATAIN_tb = 12'b0101_1000_1001;
        #10000 Rst_tb = 1;
        #11100 Rst_tb = 0;
    end
endmodule
